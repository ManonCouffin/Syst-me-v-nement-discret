-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition
-- Created on Tue Nov 30 11:39:18 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY MAEtp2 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        H : IN STD_LOGIC := '0';
        D : IN STD_LOGIC := '0';
        B : IN STD_LOGIC := '0';
        G : IN STD_LOGIC := '0';
        murD : OUT STD_LOGIC;
        murG : OUT STD_LOGIC;
        murH : OUT STD_LOGIC;
        murB : OUT STD_LOGIC
    );
END MAEtp2;

ARCHITECTURE BEHAVIOR OF MAEtp2 IS
    TYPE type_fstate IS (state2,state3,state5,state8,state9,state11,state14,state12,state1,state10,state15,state13,state16);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,H,D,B,G)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            murD <= '0';
            murG <= '0';
            murH <= '0';
            murB <= '0';
        ELSE
            murD <= '0';
            murG <= '0';
            murH <= '0';
            murB <= '0';
            CASE fstate IS
                WHEN state2 =>
                    IF (((((D = '1') AND NOT((B = '1'))) AND NOT((H = '1'))) AND NOT((G = '1')))) THEN
                        reg_fstate <= state14;
                    ELSIF ((((NOT((D = '1')) AND NOT((B = '1'))) AND (H = '1')) AND NOT((G = '1')))) THEN
                        reg_fstate <= state12;
                    ELSIF ((((NOT((D = '1')) AND (B = '1')) AND NOT((H = '1'))) AND NOT((G = '1')))) THEN
                        reg_fstate <= state8;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    murG <= '1';

                    murB <= '0';

                    murH <= '0';

                    murD <= '0';
                WHEN state3 =>
                    IF (((((B = '1') AND NOT((D = '1'))) AND NOT((G = '1'))) AND NOT((H = '1')))) THEN
                        reg_fstate <= state5;
                    ELSIF (((((D = '1') AND NOT((B = '1'))) AND NOT((H = '1'))) AND NOT((G = '1')))) THEN
                        reg_fstate <= state9;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    murG <= '1';

                    murB <= '0';

                    murH <= '1';

                    murD <= '0';
                WHEN state5 =>
                    IF (((((H = '1') AND NOT((D = '1'))) AND NOT((G = '1'))) AND NOT((B = '1')))) THEN
                        reg_fstate <= state3;
                    ELSIF (((((D = '1') AND NOT((B = '1'))) AND NOT((H = '1'))) AND NOT((G = '1')))) THEN
                        reg_fstate <= state15;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;

                    murG <= '1';

                    murB <= '1';

                    murH <= '0';

                    murD <= '0';
                WHEN state8 =>
                    IF (((((D = '1') AND NOT((B = '1'))) AND NOT((H = '1'))) AND NOT((G = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF ((((NOT((D = '1')) AND NOT((B = '1'))) AND (H = '1')) AND NOT((G = '1')))) THEN
                        reg_fstate <= state12;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state8;
                    END IF;

                    murG <= '1';

                    murB <= '1';

                    murH <= '0';

                    murD <= '0';
                WHEN state9 =>
                    IF ((((NOT((D = '1')) AND NOT((B = '1'))) AND NOT((H = '1'))) AND (G = '1'))) THEN
                        reg_fstate <= state3;
                    ELSIF ((((NOT((D = '1')) AND (B = '1')) AND NOT((H = '1'))) AND NOT((G = '1')))) THEN
                        reg_fstate <= state10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state9;
                    END IF;

                    murG <= '0';

                    murB <= '0';

                    murH <= '1';

                    murD <= '1';
                WHEN state11 =>
                    IF (((((G = '1') AND NOT((D = '1'))) AND NOT((H = '1'))) AND NOT((B = '1')))) THEN
                        reg_fstate <= state5;
                    ELSIF ((((NOT((D = '1')) AND (B = '1')) AND NOT((H = '1'))) AND NOT((G = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF (((((D = '1') AND NOT((B = '1'))) AND NOT((H = '1'))) AND NOT((G = '1')))) THEN
                        reg_fstate <= state15;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state11;
                    END IF;

                    murG <= '0';

                    murB <= '0';

                    murH <= '1';

                    murD <= '0';
                WHEN state14 =>
                    IF ((((NOT((D = '1')) AND NOT((B = '1'))) AND (H = '1')) AND NOT((G = '1')))) THEN
                        reg_fstate <= state13;
                    ELSIF ((((NOT((D = '1')) AND NOT((B = '1'))) AND NOT((H = '1'))) AND (G = '1'))) THEN
                        reg_fstate <= state2;
                    ELSIF ((((NOT((D = '1')) AND (B = '1')) AND NOT((H = '1'))) AND NOT((G = '1')))) THEN
                        reg_fstate <= state16;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state14;
                    END IF;

                    murG <= '0';

                    murB <= '0';

                    murH <= '0';

                    murD <= '1';
                WHEN state12 =>
                    IF ((((NOT((D = '1')) AND (B = '1')) AND NOT((H = '1'))) AND NOT((G = '1')))) THEN
                        reg_fstate <= state8;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state12;
                    END IF;

                    murG <= '1';

                    murB <= '0';

                    murH <= '1';

                    murD <= '1';
                WHEN state1 =>
                    IF ((((NOT((D = '1')) AND NOT((B = '1'))) AND (H = '1')) AND NOT((G = '1')))) THEN
                        reg_fstate <= state11;
                    ELSIF ((((NOT((D = '1')) AND NOT((B = '1'))) AND NOT((H = '1'))) AND (G = '1'))) THEN
                        reg_fstate <= state8;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    murG <= '0';

                    murB <= '1';

                    murH <= '0';

                    murD <= '1';
                WHEN state10 =>
                    IF ((((NOT((D = '1')) AND NOT((B = '1'))) AND (H = '1')) AND NOT((G = '1')))) THEN
                        reg_fstate <= state9;
                    ELSIF (((((D = '1') AND NOT((B = '1'))) AND NOT((H = '1'))) AND NOT((G = '1')))) THEN
                        reg_fstate <= state14;
                    ELSIF ((((NOT((D = '1')) AND NOT((B = '1'))) AND NOT((H = '1'))) AND (G = '1'))) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state10;
                    END IF;

                    murG <= '0';

                    murB <= '1';

                    murH <= '0';

                    murD <= '0';
                WHEN state15 =>
                    IF ((((NOT((D = '1')) AND NOT((B = '1'))) AND NOT((H = '1'))) AND (G = '1'))) THEN
                        reg_fstate <= state5;
                    ELSIF ((((NOT((D = '1')) AND NOT((B = '1'))) AND (H = '1')) AND NOT((G = '1')))) THEN
                        reg_fstate <= state13;
                    ELSIF ((((NOT((D = '1')) AND (B = '1')) AND NOT((H = '1'))) AND NOT((G = '1')))) THEN
                        reg_fstate <= state16;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state15;
                    END IF;

                    murG <= '0';

                    murB <= '0';

                    murH <= '0';

                    murD <= '1';
                WHEN state13 =>
                    IF ((((NOT((D = '1')) AND (B = '1')) AND NOT((H = '1'))) AND NOT((G = '1')))) THEN
                        reg_fstate <= state16;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state13;
                    END IF;

                    murG <= '1';

                    murB <= '0';

                    murH <= '1';

                    murD <= '1';
                WHEN state16 =>
                    IF ((((NOT((D = '1')) AND NOT((B = '1'))) AND (H = '1')) AND NOT((G = '1')))) THEN
                        reg_fstate <= state13;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state16;
                    END IF;

                    murG <= '1';

                    murB <= '0';

                    murH <= '1';

                    murD <= '1';
                WHEN OTHERS => 
                    murD <= 'X';
                    murG <= 'X';
                    murH <= 'X';
                    murB <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
